module bit_not (in, out);
  input in;
  wire in;
  output out;
  wire out;
  
  assign out = ~in;
  
endmodule