module bit_xor (in1, in2, out);
  input in1;
  wire in1;
  input in2;
  wire in2;
  output out;
  wire out;
  
  assign out = in1 ^ in2;
  
endmodule